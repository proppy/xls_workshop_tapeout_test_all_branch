magic
tech sky130A
magscale 1 2
timestamp 1671186313
<< viali >>
rect 1777 31297 1811 31331
rect 3985 31297 4019 31331
rect 5089 31297 5123 31331
rect 7297 31297 7331 31331
rect 8401 31297 8435 31331
rect 10609 31297 10643 31331
rect 11713 31297 11747 31331
rect 14289 31297 14323 31331
rect 15025 31297 15059 31331
rect 17233 31297 17267 31331
rect 18337 31297 18371 31331
rect 20545 31297 20579 31331
rect 22017 31297 22051 31331
rect 23857 31297 23891 31331
rect 24961 31297 24995 31331
rect 27169 31297 27203 31331
rect 28181 31297 28215 31331
rect 2421 31229 2455 31263
rect 27721 30889 27755 30923
rect 28365 30889 28399 30923
rect 1593 30685 1627 30719
rect 28365 30005 28399 30039
rect 1593 29597 1627 29631
rect 28365 29597 28399 29631
rect 1593 28509 1627 28543
rect 1593 27829 1627 27863
rect 28365 27829 28399 27863
rect 28365 27421 28399 27455
rect 1593 26333 1627 26367
rect 28365 25721 28399 25755
rect 1593 25653 1627 25687
rect 28365 25381 28399 25415
rect 1593 24157 1627 24191
rect 28365 24157 28399 24191
rect 1593 23477 1627 23511
rect 28365 23069 28399 23103
rect 1593 22389 1627 22423
rect 28365 21981 28399 22015
rect 1593 21437 1627 21471
rect 28365 21301 28399 21335
rect 1593 20213 1627 20247
rect 28365 19941 28399 19975
rect 1593 19805 1627 19839
rect 28365 19125 28399 19159
rect 1593 18037 1627 18071
rect 1593 17629 1627 17663
rect 28365 17629 28399 17663
rect 28365 16949 28399 16983
rect 1593 15997 1627 16031
rect 28365 15861 28399 15895
rect 1593 15453 1627 15487
rect 28365 14841 28399 14875
rect 1593 14365 1627 14399
rect 28365 13685 28399 13719
rect 1593 13277 1627 13311
rect 28365 13277 28399 13311
rect 1593 12189 1627 12223
rect 1593 11509 1627 11543
rect 28365 11509 28399 11543
rect 28365 11101 28399 11135
rect 1593 10013 1627 10047
rect 28365 9401 28399 9435
rect 1593 9333 1627 9367
rect 28365 9061 28399 9095
rect 1593 7837 1627 7871
rect 28365 7837 28399 7871
rect 1593 7157 1627 7191
rect 28365 6749 28399 6783
rect 1593 6069 1627 6103
rect 28365 5661 28399 5695
rect 1593 5117 1627 5151
rect 28365 4981 28399 5015
rect 1593 3893 1627 3927
rect 28365 3621 28399 3655
rect 1593 3485 1627 3519
rect 28365 2805 28399 2839
<< metal1 >>
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 1670 31288 1676 31340
rect 1728 31328 1734 31340
rect 1765 31331 1823 31337
rect 1765 31328 1777 31331
rect 1728 31300 1777 31328
rect 1728 31288 1734 31300
rect 1765 31297 1777 31300
rect 1811 31297 1823 31331
rect 1765 31291 1823 31297
rect 3878 31288 3884 31340
rect 3936 31328 3942 31340
rect 3973 31331 4031 31337
rect 3973 31328 3985 31331
rect 3936 31300 3985 31328
rect 3936 31288 3942 31300
rect 3973 31297 3985 31300
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 4982 31288 4988 31340
rect 5040 31328 5046 31340
rect 5077 31331 5135 31337
rect 5077 31328 5089 31331
rect 5040 31300 5089 31328
rect 5040 31288 5046 31300
rect 5077 31297 5089 31300
rect 5123 31297 5135 31331
rect 5077 31291 5135 31297
rect 7190 31288 7196 31340
rect 7248 31328 7254 31340
rect 7285 31331 7343 31337
rect 7285 31328 7297 31331
rect 7248 31300 7297 31328
rect 7248 31288 7254 31300
rect 7285 31297 7297 31300
rect 7331 31297 7343 31331
rect 7285 31291 7343 31297
rect 8294 31288 8300 31340
rect 8352 31328 8358 31340
rect 8389 31331 8447 31337
rect 8389 31328 8401 31331
rect 8352 31300 8401 31328
rect 8352 31288 8358 31300
rect 8389 31297 8401 31300
rect 8435 31297 8447 31331
rect 8389 31291 8447 31297
rect 10502 31288 10508 31340
rect 10560 31328 10566 31340
rect 10597 31331 10655 31337
rect 10597 31328 10609 31331
rect 10560 31300 10609 31328
rect 10560 31288 10566 31300
rect 10597 31297 10609 31300
rect 10643 31297 10655 31331
rect 10597 31291 10655 31297
rect 11606 31288 11612 31340
rect 11664 31328 11670 31340
rect 11701 31331 11759 31337
rect 11701 31328 11713 31331
rect 11664 31300 11713 31328
rect 11664 31288 11670 31300
rect 11701 31297 11713 31300
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 13814 31288 13820 31340
rect 13872 31328 13878 31340
rect 14277 31331 14335 31337
rect 14277 31328 14289 31331
rect 13872 31300 14289 31328
rect 13872 31288 13878 31300
rect 14277 31297 14289 31300
rect 14323 31297 14335 31331
rect 14277 31291 14335 31297
rect 14734 31288 14740 31340
rect 14792 31328 14798 31340
rect 15013 31331 15071 31337
rect 15013 31328 15025 31331
rect 14792 31300 15025 31328
rect 14792 31288 14798 31300
rect 15013 31297 15025 31300
rect 15059 31297 15071 31331
rect 15013 31291 15071 31297
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17221 31331 17279 31337
rect 17221 31328 17233 31331
rect 17184 31300 17233 31328
rect 17184 31288 17190 31300
rect 17221 31297 17233 31300
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 18230 31288 18236 31340
rect 18288 31328 18294 31340
rect 18325 31331 18383 31337
rect 18325 31328 18337 31331
rect 18288 31300 18337 31328
rect 18288 31288 18294 31300
rect 18325 31297 18337 31300
rect 18371 31297 18383 31331
rect 18325 31291 18383 31297
rect 20438 31288 20444 31340
rect 20496 31328 20502 31340
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 20496 31300 20545 31328
rect 20496 31288 20502 31300
rect 20533 31297 20545 31300
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 21542 31288 21548 31340
rect 21600 31328 21606 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21600 31300 22017 31328
rect 21600 31288 21606 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 23750 31288 23756 31340
rect 23808 31328 23814 31340
rect 23845 31331 23903 31337
rect 23845 31328 23857 31331
rect 23808 31300 23857 31328
rect 23808 31288 23814 31300
rect 23845 31297 23857 31300
rect 23891 31297 23903 31331
rect 23845 31291 23903 31297
rect 24854 31288 24860 31340
rect 24912 31328 24918 31340
rect 24949 31331 25007 31337
rect 24949 31328 24961 31331
rect 24912 31300 24961 31328
rect 24912 31288 24918 31300
rect 24949 31297 24961 31300
rect 24995 31297 25007 31331
rect 24949 31291 25007 31297
rect 27062 31288 27068 31340
rect 27120 31328 27126 31340
rect 27157 31331 27215 31337
rect 27157 31328 27169 31331
rect 27120 31300 27169 31328
rect 27120 31288 27126 31300
rect 27157 31297 27169 31300
rect 27203 31297 27215 31331
rect 28166 31328 28172 31340
rect 28127 31300 28172 31328
rect 27157 31291 27215 31297
rect 28166 31288 28172 31300
rect 28224 31288 28230 31340
rect 566 31220 572 31272
rect 624 31260 630 31272
rect 2409 31263 2467 31269
rect 2409 31260 2421 31263
rect 624 31232 2421 31260
rect 624 31220 630 31232
rect 2409 31229 2421 31232
rect 2455 31229 2467 31263
rect 2409 31223 2467 31229
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 27706 30920 27712 30932
rect 27667 30892 27712 30920
rect 27706 30880 27712 30892
rect 27764 30880 27770 30932
rect 28350 30920 28356 30932
rect 28311 30892 28356 30920
rect 28350 30880 28356 30892
rect 28408 30880 28414 30932
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 28350 30036 28356 30048
rect 28311 30008 28356 30036
rect 28350 29996 28356 30008
rect 28408 29996 28414 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 28350 29628 28356 29640
rect 28311 29600 28356 29628
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 28350 27860 28356 27872
rect 28311 27832 28356 27860
rect 28350 27820 28356 27832
rect 28408 27820 28414 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 28350 27452 28356 27464
rect 28311 27424 28356 27452
rect 28350 27412 28356 27424
rect 28408 27412 28414 27464
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 28350 25752 28356 25764
rect 28311 25724 28356 25752
rect 28350 25712 28356 25724
rect 28408 25712 28414 25764
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 28350 25412 28356 25424
rect 28311 25384 28356 25412
rect 28350 25372 28356 25384
rect 28408 25372 28414 25424
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 28350 24188 28356 24200
rect 28311 24160 28356 24188
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 28350 23100 28356 23112
rect 28311 23072 28356 23100
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 28350 22012 28356 22024
rect 28311 21984 28356 22012
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 1578 21468 1584 21480
rect 1539 21440 1584 21468
rect 1578 21428 1584 21440
rect 1636 21428 1642 21480
rect 28350 21332 28356 21344
rect 28311 21304 28356 21332
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 28350 19972 28356 19984
rect 28311 19944 28356 19972
rect 28350 19932 28356 19944
rect 28408 19932 28414 19984
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 28350 19156 28356 19168
rect 28311 19128 28356 19156
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 28350 16980 28356 16992
rect 28311 16952 28356 16980
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 28350 14872 28356 14884
rect 28311 14844 28356 14872
rect 28350 14832 28356 14844
rect 28408 14832 28414 14884
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 28350 13716 28356 13728
rect 28311 13688 28356 13716
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 28350 11540 28356 11552
rect 28311 11512 28356 11540
rect 28350 11500 28356 11512
rect 28408 11500 28414 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 28350 11132 28356 11144
rect 28311 11104 28356 11132
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 28350 9432 28356 9444
rect 28311 9404 28356 9432
rect 28350 9392 28356 9404
rect 28408 9392 28414 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 28350 9092 28356 9104
rect 28311 9064 28356 9092
rect 28350 9052 28356 9064
rect 28408 9052 28414 9104
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 28350 7868 28356 7880
rect 28311 7840 28356 7868
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 28350 6780 28356 6792
rect 28311 6752 28356 6780
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 28350 5692 28356 5704
rect 28311 5664 28356 5692
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 28350 5012 28356 5024
rect 28311 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 28350 3652 28356 3664
rect 28311 3624 28356 3652
rect 28350 3612 28356 3624
rect 28408 3612 28414 3664
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
<< via1 >>
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 1676 31288 1728 31340
rect 3884 31288 3936 31340
rect 4988 31288 5040 31340
rect 7196 31288 7248 31340
rect 8300 31288 8352 31340
rect 10508 31288 10560 31340
rect 11612 31288 11664 31340
rect 13820 31288 13872 31340
rect 14740 31288 14792 31340
rect 17132 31288 17184 31340
rect 18236 31288 18288 31340
rect 20444 31288 20496 31340
rect 21548 31288 21600 31340
rect 23756 31288 23808 31340
rect 24860 31288 24912 31340
rect 27068 31288 27120 31340
rect 28172 31331 28224 31340
rect 28172 31297 28181 31331
rect 28181 31297 28215 31331
rect 28215 31297 28224 31331
rect 28172 31288 28224 31297
rect 572 31220 624 31272
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 27712 30923 27764 30932
rect 27712 30889 27721 30923
rect 27721 30889 27755 30923
rect 27755 30889 27764 30923
rect 27712 30880 27764 30889
rect 28356 30923 28408 30932
rect 28356 30889 28365 30923
rect 28365 30889 28399 30923
rect 28399 30889 28408 30923
rect 28356 30880 28408 30889
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 28356 30039 28408 30048
rect 28356 30005 28365 30039
rect 28365 30005 28399 30039
rect 28399 30005 28408 30039
rect 28356 29996 28408 30005
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 28356 27863 28408 27872
rect 28356 27829 28365 27863
rect 28365 27829 28399 27863
rect 28399 27829 28408 27863
rect 28356 27820 28408 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 28356 27455 28408 27464
rect 28356 27421 28365 27455
rect 28365 27421 28399 27455
rect 28399 27421 28408 27455
rect 28356 27412 28408 27421
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 28356 25755 28408 25764
rect 28356 25721 28365 25755
rect 28365 25721 28399 25755
rect 28399 25721 28408 25755
rect 28356 25712 28408 25721
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 28356 25415 28408 25424
rect 28356 25381 28365 25415
rect 28365 25381 28399 25415
rect 28399 25381 28408 25415
rect 28356 25372 28408 25381
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 1584 21471 1636 21480
rect 1584 21437 1593 21471
rect 1593 21437 1627 21471
rect 1627 21437 1636 21471
rect 1584 21428 1636 21437
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 28356 19975 28408 19984
rect 28356 19941 28365 19975
rect 28365 19941 28399 19975
rect 28399 19941 28408 19975
rect 28356 19932 28408 19941
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 28356 16983 28408 16992
rect 28356 16949 28365 16983
rect 28365 16949 28399 16983
rect 28399 16949 28408 16983
rect 28356 16940 28408 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 28356 14875 28408 14884
rect 28356 14841 28365 14875
rect 28365 14841 28399 14875
rect 28399 14841 28408 14875
rect 28356 14832 28408 14841
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 28356 9435 28408 9444
rect 28356 9401 28365 9435
rect 28365 9401 28399 9435
rect 28399 9401 28408 9435
rect 28356 9392 28408 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 28356 9095 28408 9104
rect 28356 9061 28365 9095
rect 28365 9061 28399 9095
rect 28399 9061 28408 9095
rect 28356 9052 28408 9061
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 28356 6783 28408 6792
rect 28356 6749 28365 6783
rect 28365 6749 28399 6783
rect 28399 6749 28408 6783
rect 28356 6740 28408 6749
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 28356 3655 28408 3664
rect 28356 3621 28365 3655
rect 28365 3621 28399 3655
rect 28399 3621 28408 3655
rect 28356 3612 28408 3621
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
<< metal2 >>
rect 570 33200 626 34000
rect 1674 33200 1730 34000
rect 2778 33200 2834 34000
rect 3882 33200 3938 34000
rect 4986 33200 5042 34000
rect 6090 33200 6146 34000
rect 7194 33200 7250 34000
rect 8298 33200 8354 34000
rect 9402 33200 9458 34000
rect 10506 33200 10562 34000
rect 11610 33200 11666 34000
rect 12714 33200 12770 34000
rect 13818 33200 13874 34000
rect 14922 33200 14978 34000
rect 16026 33200 16082 34000
rect 17130 33200 17186 34000
rect 18234 33200 18290 34000
rect 19338 33200 19394 34000
rect 20442 33200 20498 34000
rect 21546 33200 21602 34000
rect 22650 33200 22706 34000
rect 23754 33200 23810 34000
rect 24858 33200 24914 34000
rect 25962 33200 26018 34000
rect 27066 33200 27122 34000
rect 28170 33200 28226 34000
rect 29274 33200 29330 34000
rect 584 31278 612 33200
rect 1688 31346 1716 33200
rect 3896 31346 3924 33200
rect 5000 31346 5028 33200
rect 7208 31346 7236 33200
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 8312 31346 8340 33200
rect 10520 31346 10548 33200
rect 11624 31346 11652 33200
rect 13832 31346 13860 33200
rect 14936 31770 14964 33200
rect 14752 31742 14964 31770
rect 14752 31346 14780 31742
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 17144 31346 17172 33200
rect 18248 31346 18276 33200
rect 20456 31346 20484 33200
rect 21560 31346 21588 33200
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 23768 31346 23796 33200
rect 24872 31346 24900 33200
rect 27080 31346 27108 33200
rect 27710 31920 27766 31929
rect 27710 31855 27766 31864
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 11612 31340 11664 31346
rect 11612 31282 11664 31288
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 14740 31340 14792 31346
rect 14740 31282 14792 31288
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 572 31272 624 31278
rect 572 31214 624 31220
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 27724 30938 27752 31855
rect 28184 31346 28212 33200
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 28354 31240 28410 31249
rect 28354 31175 28410 31184
rect 28368 30938 28396 31175
rect 27712 30932 27764 30938
rect 27712 30874 27764 30880
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 1596 30297 1624 30670
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 1582 30288 1638 30297
rect 1582 30223 1638 30232
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 28368 29889 28396 29990
rect 28354 29880 28410 29889
rect 28354 29815 28410 29824
rect 1584 29640 1636 29646
rect 1582 29608 1584 29617
rect 28356 29640 28408 29646
rect 1636 29608 1638 29617
rect 28356 29582 28408 29588
rect 1582 29543 1638 29552
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 28368 29209 28396 29582
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28354 29200 28410 29209
rect 28354 29135 28410 29144
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1596 28257 1624 28494
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 1582 28248 1638 28257
rect 7896 28251 8204 28260
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 1582 28183 1638 28192
rect 1584 27872 1636 27878
rect 28356 27872 28408 27878
rect 1584 27814 1636 27820
rect 28354 27840 28356 27849
rect 28408 27840 28410 27849
rect 1596 27577 1624 27814
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 25261 27772 25569 27781
rect 28354 27775 28410 27784
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 1582 27568 1638 27577
rect 1582 27503 1638 27512
rect 28356 27464 28408 27470
rect 28354 27432 28356 27441
rect 28408 27432 28410 27441
rect 28354 27367 28410 27376
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26217 1624 26318
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28354 25800 28410 25809
rect 28354 25735 28356 25744
rect 28408 25735 28410 25744
rect 28356 25706 28408 25712
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25537 1624 25638
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 1582 25528 1638 25537
rect 4423 25531 4731 25540
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 1582 25463 1638 25472
rect 28356 25424 28408 25430
rect 28354 25392 28356 25401
rect 28408 25392 28410 25401
rect 28354 25327 28410 25336
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 1584 24200 1636 24206
rect 1582 24168 1584 24177
rect 28356 24200 28408 24206
rect 1636 24168 1638 24177
rect 28356 24142 28408 24148
rect 1582 24103 1638 24112
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 28368 23769 28396 24142
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28354 23760 28410 23769
rect 28354 23695 28410 23704
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 28356 23112 28408 23118
rect 28354 23080 28356 23089
rect 28408 23080 28410 23089
rect 28354 23015 28410 23024
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 28356 22024 28408 22030
rect 28354 21992 28356 22001
rect 28408 21992 28410 22001
rect 28354 21927 28410 21936
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 1584 21480 1636 21486
rect 1582 21448 1584 21457
rect 1636 21448 1638 21457
rect 1582 21383 1638 21392
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 28368 21049 28396 21286
rect 28354 21040 28410 21049
rect 28354 20975 28410 20984
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 1582 20088 1638 20097
rect 4423 20091 4731 20100
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 1582 20023 1638 20032
rect 28356 19984 28408 19990
rect 28354 19952 28356 19961
rect 28408 19952 28410 19961
rect 28354 19887 28410 19896
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19417 1624 19790
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 28368 19009 28396 19110
rect 28354 19000 28410 19009
rect 28354 18935 28410 18944
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 1584 18080 1636 18086
rect 1582 18048 1584 18057
rect 1636 18048 1638 18057
rect 1582 17983 1638 17992
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 1584 17672 1636 17678
rect 28356 17672 28408 17678
rect 1584 17614 1636 17620
rect 28354 17640 28356 17649
rect 28408 17640 28410 17649
rect 1596 17377 1624 17614
rect 28354 17575 28410 17584
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 1582 17368 1638 17377
rect 7896 17371 8204 17380
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 1582 17303 1638 17312
rect 28356 16992 28408 16998
rect 28354 16960 28356 16969
rect 28408 16960 28410 16969
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 25261 16892 25569 16901
rect 28354 16895 28410 16904
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 1584 16040 1636 16046
rect 1582 16008 1584 16017
rect 1636 16008 1638 16017
rect 1582 15943 1638 15952
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 28368 15609 28396 15846
rect 28354 15600 28410 15609
rect 28354 15535 28410 15544
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15337 1624 15438
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28354 14920 28410 14929
rect 28354 14855 28356 14864
rect 28408 14855 28410 14864
rect 28356 14826 28408 14832
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 28368 13569 28396 13670
rect 28354 13560 28410 13569
rect 28354 13495 28410 13504
rect 1584 13320 1636 13326
rect 1582 13288 1584 13297
rect 28356 13320 28408 13326
rect 1636 13288 1638 13297
rect 28356 13262 28408 13268
rect 1582 13223 1638 13232
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 28368 12889 28396 13262
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11937 1624 12174
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 1582 11928 1638 11937
rect 7896 11931 8204 11940
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 1582 11863 1638 11872
rect 1584 11552 1636 11558
rect 28356 11552 28408 11558
rect 1584 11494 1636 11500
rect 28354 11520 28356 11529
rect 28408 11520 28410 11529
rect 1596 11257 1624 11494
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 25261 11452 25569 11461
rect 28354 11455 28410 11464
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 28356 11144 28408 11150
rect 28354 11112 28356 11121
rect 28408 11112 28410 11121
rect 28354 11047 28410 11056
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9897 1624 9998
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28354 9480 28410 9489
rect 28354 9415 28356 9424
rect 28408 9415 28410 9424
rect 28356 9386 28408 9392
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 1582 9208 1638 9217
rect 4423 9211 4731 9220
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 1582 9143 1638 9152
rect 28356 9104 28408 9110
rect 28354 9072 28356 9081
rect 28408 9072 28410 9081
rect 28354 9007 28410 9016
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 1584 7880 1636 7886
rect 1582 7848 1584 7857
rect 28356 7880 28408 7886
rect 1636 7848 1638 7857
rect 28356 7822 28408 7828
rect 1582 7783 1638 7792
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 28368 7449 28396 7822
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 28354 7440 28410 7449
rect 28354 7375 28410 7384
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 28356 6792 28408 6798
rect 28354 6760 28356 6769
rect 28408 6760 28410 6769
rect 28354 6695 28410 6704
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5817 1624 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 28356 5704 28408 5710
rect 28354 5672 28356 5681
rect 28408 5672 28410 5681
rect 28354 5607 28410 5616
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 1584 5160 1636 5166
rect 1582 5128 1584 5137
rect 1636 5128 1638 5137
rect 1582 5063 1638 5072
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 28368 4729 28396 4966
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3777 1624 3878
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 1582 3768 1638 3777
rect 4423 3771 4731 3780
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 1582 3703 1638 3712
rect 28356 3664 28408 3670
rect 28354 3632 28356 3641
rect 28408 3632 28410 3641
rect 28354 3567 28410 3576
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3097 1624 3470
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 28368 2689 28396 2790
rect 28354 2680 28410 2689
rect 28354 2615 28410 2624
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
<< via2 >>
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 27710 31864 27766 31920
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28354 31184 28410 31240
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 1582 30232 1638 30288
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 28354 29824 28410 29880
rect 1582 29588 1584 29608
rect 1584 29588 1636 29608
rect 1636 29588 1638 29608
rect 1582 29552 1638 29588
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28354 29144 28410 29200
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 1582 28192 1638 28248
rect 28354 27820 28356 27840
rect 28356 27820 28408 27840
rect 28408 27820 28410 27840
rect 28354 27784 28410 27820
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 1582 27512 1638 27568
rect 28354 27412 28356 27432
rect 28356 27412 28408 27432
rect 28408 27412 28410 27432
rect 28354 27376 28410 27412
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 1582 26152 1638 26208
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28354 25764 28410 25800
rect 28354 25744 28356 25764
rect 28356 25744 28408 25764
rect 28408 25744 28410 25764
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 1582 25472 1638 25528
rect 28354 25372 28356 25392
rect 28356 25372 28408 25392
rect 28408 25372 28410 25392
rect 28354 25336 28410 25372
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 1582 24148 1584 24168
rect 1584 24148 1636 24168
rect 1636 24148 1638 24168
rect 1582 24112 1638 24148
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28354 23704 28410 23760
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 28354 23060 28356 23080
rect 28356 23060 28408 23080
rect 28408 23060 28410 23080
rect 28354 23024 28410 23060
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 1582 22072 1638 22128
rect 28354 21972 28356 21992
rect 28356 21972 28408 21992
rect 28408 21972 28410 21992
rect 28354 21936 28410 21972
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 1582 21428 1584 21448
rect 1584 21428 1636 21448
rect 1636 21428 1638 21448
rect 1582 21392 1638 21428
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 28354 20984 28410 21040
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 1582 20032 1638 20088
rect 28354 19932 28356 19952
rect 28356 19932 28408 19952
rect 28408 19932 28410 19952
rect 28354 19896 28410 19932
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 1582 19352 1638 19408
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 28354 18944 28410 19000
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 1582 18028 1584 18048
rect 1584 18028 1636 18048
rect 1636 18028 1638 18048
rect 1582 17992 1638 18028
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 28354 17620 28356 17640
rect 28356 17620 28408 17640
rect 28408 17620 28410 17640
rect 28354 17584 28410 17620
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 1582 17312 1638 17368
rect 28354 16940 28356 16960
rect 28356 16940 28408 16960
rect 28408 16940 28410 16960
rect 28354 16904 28410 16940
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 1582 15988 1584 16008
rect 1584 15988 1636 16008
rect 1636 15988 1638 16008
rect 1582 15952 1638 15988
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 28354 15544 28410 15600
rect 1582 15272 1638 15328
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28354 14884 28410 14920
rect 28354 14864 28356 14884
rect 28356 14864 28408 14884
rect 28408 14864 28410 14884
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 1582 13912 1638 13968
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 28354 13504 28410 13560
rect 1582 13268 1584 13288
rect 1584 13268 1636 13288
rect 1636 13268 1638 13288
rect 1582 13232 1638 13268
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12824 28410 12880
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 1582 11872 1638 11928
rect 28354 11500 28356 11520
rect 28356 11500 28408 11520
rect 28408 11500 28410 11520
rect 28354 11464 28410 11500
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 1582 11192 1638 11248
rect 28354 11092 28356 11112
rect 28356 11092 28408 11112
rect 28408 11092 28410 11112
rect 28354 11056 28410 11092
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 1582 9832 1638 9888
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 9444 28410 9480
rect 28354 9424 28356 9444
rect 28356 9424 28408 9444
rect 28408 9424 28410 9444
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 1582 9152 1638 9208
rect 28354 9052 28356 9072
rect 28356 9052 28408 9072
rect 28408 9052 28410 9072
rect 28354 9016 28410 9052
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 1582 7828 1584 7848
rect 1584 7828 1636 7848
rect 1636 7828 1638 7848
rect 1582 7792 1638 7828
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28354 7384 28410 7440
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 28354 6740 28356 6760
rect 28356 6740 28408 6760
rect 28408 6740 28410 6760
rect 28354 6704 28410 6740
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 1582 5752 1638 5808
rect 28354 5652 28356 5672
rect 28356 5652 28408 5672
rect 28408 5652 28410 5672
rect 28354 5616 28410 5652
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 1582 5108 1584 5128
rect 1584 5108 1636 5128
rect 1636 5108 1638 5128
rect 1582 5072 1638 5108
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 28354 4664 28410 4720
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 1582 3712 1638 3768
rect 28354 3612 28356 3632
rect 28356 3612 28408 3632
rect 28408 3612 28410 3632
rect 28354 3576 28410 3612
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 1582 3032 1638 3088
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28354 2624 28410 2680
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 27705 31922 27771 31925
rect 29200 31922 30000 31952
rect 27705 31920 30000 31922
rect 27705 31864 27710 31920
rect 27766 31864 30000 31920
rect 27705 31862 30000 31864
rect 27705 31859 27771 31862
rect 29200 31832 30000 31862
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 28349 31242 28415 31245
rect 29200 31242 30000 31272
rect 28349 31240 30000 31242
rect 28349 31184 28354 31240
rect 28410 31184 30000 31240
rect 28349 31182 30000 31184
rect 28349 31179 28415 31182
rect 29200 31152 30000 31182
rect 4419 31040 4735 31041
rect 0 30880 800 31000
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 29200 30472 30000 30592
rect 28730 30431 29046 30432
rect 0 30290 800 30320
rect 1577 30290 1643 30293
rect 0 30288 1643 30290
rect 0 30232 1582 30288
rect 1638 30232 1643 30288
rect 0 30230 1643 30232
rect 0 30200 800 30230
rect 1577 30227 1643 30230
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 28349 29882 28415 29885
rect 29200 29882 30000 29912
rect 28349 29880 30000 29882
rect 28349 29824 28354 29880
rect 28410 29824 30000 29880
rect 28349 29822 30000 29824
rect 28349 29819 28415 29822
rect 29200 29792 30000 29822
rect 0 29610 800 29640
rect 1577 29610 1643 29613
rect 0 29608 1643 29610
rect 0 29552 1582 29608
rect 1638 29552 1643 29608
rect 0 29550 1643 29552
rect 0 29520 800 29550
rect 1577 29547 1643 29550
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 28349 29202 28415 29205
rect 29200 29202 30000 29232
rect 28349 29200 30000 29202
rect 28349 29144 28354 29200
rect 28410 29144 30000 29200
rect 28349 29142 30000 29144
rect 28349 29139 28415 29142
rect 29200 29112 30000 29142
rect 0 28840 800 28960
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 29200 28432 30000 28552
rect 7892 28320 8208 28321
rect 0 28250 800 28280
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 1577 28250 1643 28253
rect 0 28248 1643 28250
rect 0 28192 1582 28248
rect 1638 28192 1643 28248
rect 0 28190 1643 28192
rect 0 28160 800 28190
rect 1577 28187 1643 28190
rect 28349 27842 28415 27845
rect 29200 27842 30000 27872
rect 28349 27840 30000 27842
rect 28349 27784 28354 27840
rect 28410 27784 30000 27840
rect 28349 27782 30000 27784
rect 28349 27779 28415 27782
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 29200 27752 30000 27782
rect 25257 27711 25573 27712
rect 0 27570 800 27600
rect 1577 27570 1643 27573
rect 0 27568 1643 27570
rect 0 27512 1582 27568
rect 1638 27512 1643 27568
rect 0 27510 1643 27512
rect 0 27480 800 27510
rect 1577 27507 1643 27510
rect 28349 27434 28415 27437
rect 28349 27432 29378 27434
rect 28349 27376 28354 27432
rect 28410 27376 29378 27432
rect 28349 27374 29378 27376
rect 28349 27371 28415 27374
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 29318 27192 29378 27374
rect 28730 27167 29046 27168
rect 29200 27072 30000 27192
rect 0 26800 800 26920
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 29200 26392 30000 26512
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 28349 25802 28415 25805
rect 29200 25802 30000 25832
rect 28349 25800 30000 25802
rect 28349 25744 28354 25800
rect 28410 25744 30000 25800
rect 28349 25742 30000 25744
rect 28349 25739 28415 25742
rect 29200 25712 30000 25742
rect 4419 25600 4735 25601
rect 0 25530 800 25560
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 1577 25530 1643 25533
rect 0 25528 1643 25530
rect 0 25472 1582 25528
rect 1638 25472 1643 25528
rect 0 25470 1643 25472
rect 0 25440 800 25470
rect 1577 25467 1643 25470
rect 28349 25394 28415 25397
rect 28349 25392 29378 25394
rect 28349 25336 28354 25392
rect 28410 25336 29378 25392
rect 28349 25334 29378 25336
rect 28349 25331 28415 25334
rect 29318 25152 29378 25334
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 29200 25032 30000 25152
rect 28730 24991 29046 24992
rect 0 24760 800 24880
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 29200 24352 30000 24472
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 28349 23762 28415 23765
rect 29200 23762 30000 23792
rect 28349 23760 30000 23762
rect 28349 23704 28354 23760
rect 28410 23704 30000 23760
rect 28349 23702 30000 23704
rect 28349 23699 28415 23702
rect 29200 23672 30000 23702
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 28349 23082 28415 23085
rect 29200 23082 30000 23112
rect 28349 23080 30000 23082
rect 28349 23024 28354 23080
rect 28410 23024 30000 23080
rect 28349 23022 30000 23024
rect 28349 23019 28415 23022
rect 29200 22992 30000 23022
rect 7892 22880 8208 22881
rect 0 22720 800 22840
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 29200 22312 30000 22432
rect 25257 22271 25573 22272
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 28349 21994 28415 21997
rect 28349 21992 29378 21994
rect 28349 21936 28354 21992
rect 28410 21936 29378 21992
rect 28349 21934 29378 21936
rect 28349 21931 28415 21934
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 29318 21752 29378 21934
rect 28730 21727 29046 21728
rect 29200 21632 30000 21752
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 0 20680 800 20800
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 29200 20272 30000 20392
rect 4419 20160 4735 20161
rect 0 20090 800 20120
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 28349 19954 28415 19957
rect 28349 19952 29378 19954
rect 28349 19896 28354 19952
rect 28410 19896 29378 19952
rect 28349 19894 29378 19896
rect 28349 19891 28415 19894
rect 29318 19712 29378 19894
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 29200 19592 30000 19712
rect 28730 19551 29046 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 28349 19002 28415 19005
rect 29200 19002 30000 19032
rect 28349 19000 30000 19002
rect 28349 18944 28354 19000
rect 28410 18944 30000 19000
rect 28349 18942 30000 18944
rect 28349 18939 28415 18942
rect 29200 18912 30000 18942
rect 0 18640 800 18760
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 29200 18232 30000 18352
rect 0 18050 800 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 800 17990
rect 1577 17987 1643 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 28349 17642 28415 17645
rect 29200 17642 30000 17672
rect 28349 17640 30000 17642
rect 28349 17584 28354 17640
rect 28410 17584 30000 17640
rect 28349 17582 30000 17584
rect 28349 17579 28415 17582
rect 29200 17552 30000 17582
rect 7892 17440 8208 17441
rect 0 17370 800 17400
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 28349 16962 28415 16965
rect 29200 16962 30000 16992
rect 28349 16960 30000 16962
rect 28349 16904 28354 16960
rect 28410 16904 30000 16960
rect 28349 16902 30000 16904
rect 28349 16899 28415 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 29200 16872 30000 16902
rect 25257 16831 25573 16832
rect 0 16600 800 16720
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 29200 16192 30000 16312
rect 0 16010 800 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 800 15950
rect 1577 15947 1643 15950
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 28349 15602 28415 15605
rect 29200 15602 30000 15632
rect 28349 15600 30000 15602
rect 28349 15544 28354 15600
rect 28410 15544 30000 15600
rect 28349 15542 30000 15544
rect 28349 15539 28415 15542
rect 29200 15512 30000 15542
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 28349 14922 28415 14925
rect 29200 14922 30000 14952
rect 28349 14920 30000 14922
rect 28349 14864 28354 14920
rect 28410 14864 30000 14920
rect 28349 14862 30000 14864
rect 28349 14859 28415 14862
rect 29200 14832 30000 14862
rect 4419 14720 4735 14721
rect 0 14560 800 14680
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 29200 14152 30000 14272
rect 28730 14111 29046 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 28349 13562 28415 13565
rect 29200 13562 30000 13592
rect 28349 13560 30000 13562
rect 28349 13504 28354 13560
rect 28410 13504 30000 13560
rect 28349 13502 30000 13504
rect 28349 13499 28415 13502
rect 29200 13472 30000 13502
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 28349 12882 28415 12885
rect 29200 12882 30000 12912
rect 28349 12880 30000 12882
rect 28349 12824 28354 12880
rect 28410 12824 30000 12880
rect 28349 12822 30000 12824
rect 28349 12819 28415 12822
rect 29200 12792 30000 12822
rect 0 12520 800 12640
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 29200 12112 30000 12232
rect 7892 12000 8208 12001
rect 0 11930 800 11960
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 800 11870
rect 1577 11867 1643 11870
rect 28349 11522 28415 11525
rect 29200 11522 30000 11552
rect 28349 11520 30000 11522
rect 28349 11464 28354 11520
rect 28410 11464 30000 11520
rect 28349 11462 30000 11464
rect 28349 11459 28415 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 29200 11432 30000 11462
rect 25257 11391 25573 11392
rect 0 11250 800 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 800 11190
rect 1577 11187 1643 11190
rect 28349 11114 28415 11117
rect 28349 11112 29378 11114
rect 28349 11056 28354 11112
rect 28410 11056 29378 11112
rect 28349 11054 29378 11056
rect 28349 11051 28415 11054
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 29318 10872 29378 11054
rect 28730 10847 29046 10848
rect 29200 10752 30000 10872
rect 0 10480 800 10600
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 29200 10072 30000 10192
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 28349 9482 28415 9485
rect 29200 9482 30000 9512
rect 28349 9480 30000 9482
rect 28349 9424 28354 9480
rect 28410 9424 30000 9480
rect 28349 9422 30000 9424
rect 28349 9419 28415 9422
rect 29200 9392 30000 9422
rect 4419 9280 4735 9281
rect 0 9210 800 9240
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 28349 9074 28415 9077
rect 28349 9072 29378 9074
rect 28349 9016 28354 9072
rect 28410 9016 29378 9072
rect 28349 9014 29378 9016
rect 28349 9011 28415 9014
rect 29318 8832 29378 9014
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 29200 8712 30000 8832
rect 28730 8671 29046 8672
rect 0 8440 800 8560
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 29200 8032 30000 8152
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 28349 7442 28415 7445
rect 29200 7442 30000 7472
rect 28349 7440 30000 7442
rect 28349 7384 28354 7440
rect 28410 7384 30000 7440
rect 28349 7382 30000 7384
rect 28349 7379 28415 7382
rect 29200 7352 30000 7382
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 28349 6762 28415 6765
rect 29200 6762 30000 6792
rect 28349 6760 30000 6762
rect 28349 6704 28354 6760
rect 28410 6704 30000 6760
rect 28349 6702 30000 6704
rect 28349 6699 28415 6702
rect 29200 6672 30000 6702
rect 7892 6560 8208 6561
rect 0 6400 800 6520
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 29200 5992 30000 6112
rect 25257 5951 25573 5952
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 28349 5674 28415 5677
rect 28349 5672 29378 5674
rect 28349 5616 28354 5672
rect 28410 5616 29378 5672
rect 28349 5614 29378 5616
rect 28349 5611 28415 5614
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 29318 5432 29378 5614
rect 28730 5407 29046 5408
rect 29200 5312 30000 5432
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 28349 4722 28415 4725
rect 29200 4722 30000 4752
rect 28349 4720 30000 4722
rect 28349 4664 28354 4720
rect 28410 4664 30000 4720
rect 28349 4662 30000 4664
rect 28349 4659 28415 4662
rect 29200 4632 30000 4662
rect 0 4360 800 4480
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 29200 3952 30000 4072
rect 4419 3840 4735 3841
rect 0 3770 800 3800
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 28349 3634 28415 3637
rect 28349 3632 29378 3634
rect 28349 3576 28354 3632
rect 28410 3576 29378 3632
rect 28349 3574 29378 3576
rect 28349 3571 28415 3574
rect 29318 3392 29378 3574
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 29200 3272 30000 3392
rect 28730 3231 29046 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 28349 2682 28415 2685
rect 29200 2682 30000 2712
rect 28349 2680 30000 2682
rect 28349 2624 28354 2680
rect 28410 2624 30000 2680
rect 28349 2622 30000 2624
rect 28349 2619 28415 2622
rect 29200 2592 30000 2622
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 29200 1912 30000 2032
<< via3 >>
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 31040 4737 31600
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 31584 8210 31600
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 31040 11683 31600
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 31584 15156 31600
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 31040 18629 31600
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 31584 22102 31600
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 31040 25575 31600
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 31584 29048 31600
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1666464484
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1666464484
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_293
timestamp 1666464484
transform 1 0 28060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1666464484
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1666464484
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1666464484
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_293
timestamp 1666464484
transform 1 0 28060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1666464484
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1666464484
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1666464484
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1666464484
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1666464484
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1666464484
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1666464484
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1666464484
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1666464484
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1666464484
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1666464484
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1666464484
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1666464484
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1666464484
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_8
timestamp 1666464484
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1666464484
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1666464484
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666464484
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666464484
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666464484
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_289
timestamp 1666464484
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1666464484
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_293
timestamp 1666464484
transform 1 0 28060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1666464484
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1666464484
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_293
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1666464484
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1666464484
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1666464484
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1666464484
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666464484
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_293
timestamp 1666464484
transform 1 0 28060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666464484
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1666464484
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_293
timestamp 1666464484
transform 1 0 28060 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1666464484
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1666464484
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1666464484
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1666464484
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666464484
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666464484
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666464484
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1666464484
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1666464484
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1666464484
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1666464484
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_32
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1666464484
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1666464484
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1666464484
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1666464484
transform 1 0 28060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1666464484
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_8
timestamp 1666464484
transform 1 0 1840 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_20
timestamp 1666464484
transform 1 0 2944 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_32
timestamp 1666464484
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1666464484
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1666464484
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1666464484
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1666464484
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_293
timestamp 1666464484
transform 1 0 28060 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1666464484
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1666464484
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1666464484
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1666464484
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1666464484
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1666464484
transform 1 0 28428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_8
timestamp 1666464484
transform 1 0 1840 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1666464484
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1666464484
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1666464484
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1666464484
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_293
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1666464484
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1666464484
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1666464484
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1666464484
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_285
timestamp 1666464484
transform 1 0 27324 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1666464484
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1666464484
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_10
timestamp 1666464484
transform 1 0 2024 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_17
timestamp 1666464484
transform 1 0 2668 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_25
timestamp 1666464484
transform 1 0 3404 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_29
timestamp 1666464484
transform 1 0 3772 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_34
timestamp 1666464484
transform 1 0 4232 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_42
timestamp 1666464484
transform 1 0 4968 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_46
timestamp 1666464484
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1666464484
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_65
timestamp 1666464484
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_70
timestamp 1666464484
transform 1 0 7544 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_78
timestamp 1666464484
transform 1 0 8280 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_82
timestamp 1666464484
transform 1 0 8648 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_85
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_97
timestamp 1666464484
transform 1 0 10028 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_106
timestamp 1666464484
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_118
timestamp 1666464484
transform 1 0 11960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_130
timestamp 1666464484
transform 1 0 13064 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_138
timestamp 1666464484
transform 1 0 13800 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_141
timestamp 1666464484
transform 1 0 14076 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_146
timestamp 1666464484
transform 1 0 14536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_150
timestamp 1666464484
transform 1 0 14904 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_154
timestamp 1666464484
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_178
timestamp 1666464484
transform 1 0 17480 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_186
timestamp 1666464484
transform 1 0 18216 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_190
timestamp 1666464484
transform 1 0 18584 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_197
timestamp 1666464484
transform 1 0 19228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1666464484
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1666464484
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1666464484
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_230
timestamp 1666464484
transform 1 0 22264 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_242
timestamp 1666464484
transform 1 0 23368 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_250
timestamp 1666464484
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_262
timestamp 1666464484
transform 1 0 25208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1666464484
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_286
timestamp 1666464484
transform 1 0 27416 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 3680 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 13984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_2
timestamp 1666464484
transform 1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_3
timestamp 1666464484
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_4
timestamp 1666464484
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_5
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_6
timestamp 1666464484
transform 1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_7
timestamp 1666464484
transform 1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_8
timestamp 1666464484
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_9
timestamp 1666464484
transform 1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_10
timestamp 1666464484
transform 1 0 28152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_11
timestamp 1666464484
transform 1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_12
timestamp 1666464484
transform 1 0 28152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_13
timestamp 1666464484
transform 1 0 28152 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_14
timestamp 1666464484
transform -1 0 28428 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_15
timestamp 1666464484
transform -1 0 25208 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_16
timestamp 1666464484
transform -1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_17
timestamp 1666464484
transform -1 0 18584 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_18
timestamp 1666464484
transform -1 0 15272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_19
timestamp 1666464484
transform -1 0 11960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_20
timestamp 1666464484
transform -1 0 8648 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_21
timestamp 1666464484
transform -1 0 5336 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_22
timestamp 1666464484
transform -1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_23
timestamp 1666464484
transform -1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24
timestamp 1666464484
transform -1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform -1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform -1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform -1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform 1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform 1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform 1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform 1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform 1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform 1 0 28152 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform 1 0 27508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform -1 0 27416 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform -1 0 24104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform -1 0 20792 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform -1 0 17480 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform -1 0 14536 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform -1 0 7544 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform -1 0 4232 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform -1 0 2668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform -1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform -1 0 1840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform -1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform 1 0 28152 0 -1 5440
box -38 -48 314 592
<< labels >>
flabel metal3 s 29200 1912 30000 2032 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 29200 22312 30000 22432 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 29200 24352 30000 24472 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 29200 26392 30000 26512 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 29200 28432 30000 28552 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 29200 30472 30000 30592 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 29274 33200 29330 34000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 25962 33200 26018 34000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 22650 33200 22706 34000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 19338 33200 19394 34000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 16026 33200 16082 34000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 29200 3952 30000 4072 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 12714 33200 12770 34000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 9402 33200 9458 34000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 6090 33200 6146 34000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 2778 33200 2834 34000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 29200 5992 30000 6112 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 29200 8032 30000 8152 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 29200 10072 30000 10192 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 29200 12112 30000 12232 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 29200 14152 30000 14272 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 29200 16192 30000 16312 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 29200 18232 30000 18352 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 29200 20272 30000 20392 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 29200 3272 30000 3392 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 29200 23672 30000 23792 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 29200 25712 30000 25832 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 29200 27752 30000 27872 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 29200 29792 30000 29912 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 29200 31832 30000 31952 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 27066 33200 27122 34000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 23754 33200 23810 34000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 20442 33200 20498 34000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 17130 33200 17186 34000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 13818 33200 13874 34000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 29200 5312 30000 5432 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 10506 33200 10562 34000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 7194 33200 7250 34000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 3882 33200 3938 34000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 570 33200 626 34000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 29200 9392 30000 9512 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 29200 11432 30000 11552 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 29200 13472 30000 13592 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 29200 15512 30000 15632 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 29200 17552 30000 17672 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 29200 19592 30000 19712 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 29200 21632 30000 21752 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 29200 2592 30000 2712 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 29200 22992 30000 23112 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 29200 25032 30000 25152 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 29200 27072 30000 27192 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 29200 29112 30000 29232 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 29200 31152 30000 31272 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 28170 33200 28226 34000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 24858 33200 24914 34000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 21546 33200 21602 34000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 18234 33200 18290 34000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 14922 33200 14978 34000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 29200 4632 30000 4752 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 11610 33200 11666 34000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 8298 33200 8354 34000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 4986 33200 5042 34000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 1674 33200 1730 34000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 29200 6672 30000 6792 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 29200 10752 30000 10872 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 29200 12792 30000 12912 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 29200 14832 30000 14952 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 29200 16872 30000 16992 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 29200 18912 30000 19032 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4417 2128 4737 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 11363 2128 11683 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 18309 2128 18629 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 25255 2128 25575 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7890 2128 8210 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 14996 31008 14996 31008 0 vccd1
rlabel via1 15076 31552 15076 31552 0 vssd1
rlabel via2 28382 6749 28382 6749 0 net1
rlabel via2 28382 25381 28382 25381 0 net10
rlabel via2 28382 27421 28382 27421 0 net11
rlabel metal2 28382 29393 28382 29393 0 net12
rlabel metal2 28382 31059 28382 31059 0 net13
rlabel metal2 28198 32276 28198 32276 0 net14
rlabel metal1 24932 31314 24932 31314 0 net15
rlabel metal1 21804 31314 21804 31314 0 net16
rlabel metal1 18308 31314 18308 31314 0 net17
rlabel metal1 14904 31314 14904 31314 0 net18
rlabel metal1 11684 31314 11684 31314 0 net19
rlabel via2 28382 9061 28382 9061 0 net2
rlabel metal1 8372 31314 8372 31314 0 net20
rlabel metal1 5060 31314 5060 31314 0 net21
rlabel metal1 1748 31314 1748 31314 0 net22
rlabel metal3 1142 30260 1142 30260 0 net23
rlabel metal3 1142 28220 1142 28220 0 net24
rlabel metal3 1142 26180 1142 26180 0 net25
rlabel metal3 1142 24140 1142 24140 0 net26
rlabel metal3 1142 22100 1142 22100 0 net27
rlabel metal3 1142 20060 1142 20060 0 net28
rlabel metal3 1142 18020 1142 18020 0 net29
rlabel via2 28382 11101 28382 11101 0 net3
rlabel metal3 1142 15980 1142 15980 0 net30
rlabel metal3 1142 13940 1142 13940 0 net31
rlabel metal3 1142 11900 1142 11900 0 net32
rlabel metal3 1142 9860 1142 9860 0 net33
rlabel metal3 1142 7820 1142 7820 0 net34
rlabel metal3 1142 5780 1142 5780 0 net35
rlabel metal3 1142 3740 1142 3740 0 net36
rlabel via2 28382 3621 28382 3621 0 net37
rlabel via2 28382 5661 28382 5661 0 net38
rlabel metal2 28382 7633 28382 7633 0 net39
rlabel metal2 28382 13073 28382 13073 0 net4
rlabel via2 28382 9435 28382 9435 0 net40
rlabel via2 28382 11509 28382 11509 0 net41
rlabel metal2 28382 13617 28382 13617 0 net42
rlabel metal2 28382 15725 28382 15725 0 net43
rlabel via2 28382 17629 28382 17629 0 net44
rlabel via2 28382 19941 28382 19941 0 net45
rlabel via2 28382 21981 28382 21981 0 net46
rlabel metal2 28382 23953 28382 23953 0 net47
rlabel via2 28382 25755 28382 25755 0 net48
rlabel via2 28382 27829 28382 27829 0 net49
rlabel via2 28382 14875 28382 14875 0 net5
rlabel metal2 28382 29937 28382 29937 0 net50
rlabel metal3 28528 31892 28528 31892 0 net51
rlabel metal1 27140 31314 27140 31314 0 net52
rlabel metal1 23828 31314 23828 31314 0 net53
rlabel metal1 20516 31314 20516 31314 0 net54
rlabel metal1 17204 31314 17204 31314 0 net55
rlabel metal1 14076 31314 14076 31314 0 net56
rlabel metal1 10580 31314 10580 31314 0 net57
rlabel metal1 7268 31314 7268 31314 0 net58
rlabel metal1 3956 31314 3956 31314 0 net59
rlabel via2 28382 16949 28382 16949 0 net6
rlabel metal1 1518 31246 1518 31246 0 net60
rlabel metal3 1142 29580 1142 29580 0 net61
rlabel metal3 1142 27540 1142 27540 0 net62
rlabel metal3 1142 25500 1142 25500 0 net63
rlabel metal3 1142 23460 1142 23460 0 net64
rlabel metal3 1142 21420 1142 21420 0 net65
rlabel metal3 1142 19380 1142 19380 0 net66
rlabel metal3 1142 17340 1142 17340 0 net67
rlabel metal3 1142 15300 1142 15300 0 net68
rlabel metal3 1142 13260 1142 13260 0 net69
rlabel metal2 28382 19057 28382 19057 0 net7
rlabel metal3 1142 11220 1142 11220 0 net70
rlabel metal3 1142 9180 1142 9180 0 net71
rlabel metal3 1142 7140 1142 7140 0 net72
rlabel metal3 1142 5100 1142 5100 0 net73
rlabel metal3 1142 3060 1142 3060 0 net74
rlabel metal3 28850 2652 28850 2652 0 net75
rlabel metal2 28382 4845 28382 4845 0 net76
rlabel metal2 28382 21165 28382 21165 0 net8
rlabel via2 28382 23069 28382 23069 0 net9
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>
