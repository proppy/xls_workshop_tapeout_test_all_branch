magic
tech sky130A
magscale 1 2
timestamp 1671184448
<< nwell >>
rect 1066 30725 28926 31291
rect 1066 29637 28926 30203
rect 1066 28549 28926 29115
rect 1066 27461 28926 28027
rect 1066 26373 28926 26939
rect 1066 25285 28926 25851
rect 1066 24197 28926 24763
rect 1066 23109 28926 23675
rect 1066 22021 28926 22587
rect 1066 20933 28926 21499
rect 1066 19845 28926 20411
rect 1066 18757 28926 19323
rect 1066 17669 28926 18235
rect 1066 16581 28926 17147
rect 1066 15493 28926 16059
rect 1066 14405 28926 14971
rect 1066 13317 28926 13883
rect 1066 12229 28926 12795
rect 1066 11141 28926 11707
rect 1066 10053 28926 10619
rect 1066 8965 28926 9531
rect 1066 7877 28926 8443
rect 1066 6789 28926 7355
rect 1066 5701 28926 6267
rect 1066 4613 28926 5179
rect 1066 3525 28926 4091
rect 1066 2437 28926 3003
<< obsli1 >>
rect 1104 2159 28888 31569
<< obsm1 >>
rect 1104 2128 29048 31884
<< metal2 >>
rect 4526 33200 4582 34000
rect 4710 33200 4766 34000
rect 4894 33200 4950 34000
rect 5078 33200 5134 34000
rect 5262 33200 5318 34000
rect 5446 33200 5502 34000
rect 5630 33200 5686 34000
rect 5814 33200 5870 34000
rect 5998 33200 6054 34000
rect 6182 33200 6238 34000
rect 6366 33200 6422 34000
rect 6550 33200 6606 34000
rect 6734 33200 6790 34000
rect 6918 33200 6974 34000
rect 7102 33200 7158 34000
rect 7286 33200 7342 34000
rect 7470 33200 7526 34000
rect 7654 33200 7710 34000
rect 7838 33200 7894 34000
rect 8022 33200 8078 34000
rect 8206 33200 8262 34000
rect 8390 33200 8446 34000
rect 8574 33200 8630 34000
rect 8758 33200 8814 34000
rect 8942 33200 8998 34000
rect 9126 33200 9182 34000
rect 9310 33200 9366 34000
rect 9494 33200 9550 34000
rect 9678 33200 9734 34000
rect 9862 33200 9918 34000
rect 10046 33200 10102 34000
rect 10230 33200 10286 34000
rect 10414 33200 10470 34000
rect 10598 33200 10654 34000
rect 10782 33200 10838 34000
rect 10966 33200 11022 34000
rect 11150 33200 11206 34000
rect 11334 33200 11390 34000
rect 11518 33200 11574 34000
rect 11702 33200 11758 34000
rect 11886 33200 11942 34000
rect 12070 33200 12126 34000
rect 12254 33200 12310 34000
rect 12438 33200 12494 34000
rect 12622 33200 12678 34000
rect 12806 33200 12862 34000
rect 12990 33200 13046 34000
rect 13174 33200 13230 34000
rect 13358 33200 13414 34000
rect 13542 33200 13598 34000
rect 13726 33200 13782 34000
rect 13910 33200 13966 34000
rect 14094 33200 14150 34000
rect 14278 33200 14334 34000
rect 14462 33200 14518 34000
rect 14646 33200 14702 34000
rect 14830 33200 14886 34000
rect 15014 33200 15070 34000
rect 15198 33200 15254 34000
rect 15382 33200 15438 34000
rect 15566 33200 15622 34000
rect 15750 33200 15806 34000
rect 15934 33200 15990 34000
rect 16118 33200 16174 34000
rect 16302 33200 16358 34000
rect 16486 33200 16542 34000
rect 16670 33200 16726 34000
rect 16854 33200 16910 34000
rect 17038 33200 17094 34000
rect 17222 33200 17278 34000
rect 17406 33200 17462 34000
rect 17590 33200 17646 34000
rect 17774 33200 17830 34000
rect 17958 33200 18014 34000
rect 18142 33200 18198 34000
rect 18326 33200 18382 34000
rect 18510 33200 18566 34000
rect 18694 33200 18750 34000
rect 18878 33200 18934 34000
rect 19062 33200 19118 34000
rect 19246 33200 19302 34000
rect 19430 33200 19486 34000
rect 19614 33200 19670 34000
rect 19798 33200 19854 34000
rect 19982 33200 20038 34000
rect 20166 33200 20222 34000
rect 20350 33200 20406 34000
rect 20534 33200 20590 34000
rect 20718 33200 20774 34000
rect 20902 33200 20958 34000
rect 21086 33200 21142 34000
rect 21270 33200 21326 34000
rect 21454 33200 21510 34000
rect 21638 33200 21694 34000
rect 21822 33200 21878 34000
rect 22006 33200 22062 34000
rect 22190 33200 22246 34000
rect 22374 33200 22430 34000
rect 22558 33200 22614 34000
rect 22742 33200 22798 34000
rect 22926 33200 22982 34000
rect 23110 33200 23166 34000
rect 23294 33200 23350 34000
rect 23478 33200 23534 34000
rect 23662 33200 23718 34000
rect 23846 33200 23902 34000
rect 24030 33200 24086 34000
rect 24214 33200 24270 34000
rect 24398 33200 24454 34000
rect 24582 33200 24638 34000
rect 24766 33200 24822 34000
rect 24950 33200 25006 34000
rect 25134 33200 25190 34000
rect 25318 33200 25374 34000
<< obsm2 >>
rect 4423 33144 4470 33200
rect 4638 33144 4654 33200
rect 4822 33144 4838 33200
rect 5006 33144 5022 33200
rect 5190 33144 5206 33200
rect 5374 33144 5390 33200
rect 5558 33144 5574 33200
rect 5742 33144 5758 33200
rect 5926 33144 5942 33200
rect 6110 33144 6126 33200
rect 6294 33144 6310 33200
rect 6478 33144 6494 33200
rect 6662 33144 6678 33200
rect 6846 33144 6862 33200
rect 7030 33144 7046 33200
rect 7214 33144 7230 33200
rect 7398 33144 7414 33200
rect 7582 33144 7598 33200
rect 7766 33144 7782 33200
rect 7950 33144 7966 33200
rect 8134 33144 8150 33200
rect 8318 33144 8334 33200
rect 8502 33144 8518 33200
rect 8686 33144 8702 33200
rect 8870 33144 8886 33200
rect 9054 33144 9070 33200
rect 9238 33144 9254 33200
rect 9422 33144 9438 33200
rect 9606 33144 9622 33200
rect 9790 33144 9806 33200
rect 9974 33144 9990 33200
rect 10158 33144 10174 33200
rect 10342 33144 10358 33200
rect 10526 33144 10542 33200
rect 10710 33144 10726 33200
rect 10894 33144 10910 33200
rect 11078 33144 11094 33200
rect 11262 33144 11278 33200
rect 11446 33144 11462 33200
rect 11630 33144 11646 33200
rect 11814 33144 11830 33200
rect 11998 33144 12014 33200
rect 12182 33144 12198 33200
rect 12366 33144 12382 33200
rect 12550 33144 12566 33200
rect 12734 33144 12750 33200
rect 12918 33144 12934 33200
rect 13102 33144 13118 33200
rect 13286 33144 13302 33200
rect 13470 33144 13486 33200
rect 13654 33144 13670 33200
rect 13838 33144 13854 33200
rect 14022 33144 14038 33200
rect 14206 33144 14222 33200
rect 14390 33144 14406 33200
rect 14574 33144 14590 33200
rect 14758 33144 14774 33200
rect 14942 33144 14958 33200
rect 15126 33144 15142 33200
rect 15310 33144 15326 33200
rect 15494 33144 15510 33200
rect 15678 33144 15694 33200
rect 15862 33144 15878 33200
rect 16046 33144 16062 33200
rect 16230 33144 16246 33200
rect 16414 33144 16430 33200
rect 16598 33144 16614 33200
rect 16782 33144 16798 33200
rect 16966 33144 16982 33200
rect 17150 33144 17166 33200
rect 17334 33144 17350 33200
rect 17518 33144 17534 33200
rect 17702 33144 17718 33200
rect 17886 33144 17902 33200
rect 18070 33144 18086 33200
rect 18254 33144 18270 33200
rect 18438 33144 18454 33200
rect 18622 33144 18638 33200
rect 18806 33144 18822 33200
rect 18990 33144 19006 33200
rect 19174 33144 19190 33200
rect 19358 33144 19374 33200
rect 19542 33144 19558 33200
rect 19726 33144 19742 33200
rect 19910 33144 19926 33200
rect 20094 33144 20110 33200
rect 20278 33144 20294 33200
rect 20462 33144 20478 33200
rect 20646 33144 20662 33200
rect 20830 33144 20846 33200
rect 21014 33144 21030 33200
rect 21198 33144 21214 33200
rect 21382 33144 21398 33200
rect 21566 33144 21582 33200
rect 21750 33144 21766 33200
rect 21934 33144 21950 33200
rect 22118 33144 22134 33200
rect 22302 33144 22318 33200
rect 22486 33144 22502 33200
rect 22670 33144 22686 33200
rect 22854 33144 22870 33200
rect 23038 33144 23054 33200
rect 23222 33144 23238 33200
rect 23406 33144 23422 33200
rect 23590 33144 23606 33200
rect 23774 33144 23790 33200
rect 23958 33144 23974 33200
rect 24142 33144 24158 33200
rect 24326 33144 24342 33200
rect 24510 33144 24526 33200
rect 24694 33144 24710 33200
rect 24878 33144 24894 33200
rect 25062 33144 25078 33200
rect 25246 33144 25262 33200
rect 25430 33144 29042 33200
rect 4423 2139 29042 33144
<< obsm3 >>
rect 4419 2143 29046 31585
<< metal4 >>
rect 4417 2128 4737 31600
rect 7890 2128 8210 31600
rect 11363 2128 11683 31600
rect 14836 2128 15156 31600
rect 18309 2128 18629 31600
rect 21782 2128 22102 31600
rect 25255 2128 25575 31600
rect 28728 2128 29048 31600
<< labels >>
rlabel metal2 s 4526 33200 4582 34000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 10046 33200 10102 34000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 10598 33200 10654 34000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 11150 33200 11206 34000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 11702 33200 11758 34000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 12254 33200 12310 34000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 12806 33200 12862 34000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 13358 33200 13414 34000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 13910 33200 13966 34000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 14462 33200 14518 34000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 15014 33200 15070 34000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5078 33200 5134 34000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 15566 33200 15622 34000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 16118 33200 16174 34000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 16670 33200 16726 34000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 17222 33200 17278 34000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 17774 33200 17830 34000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 18326 33200 18382 34000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 18878 33200 18934 34000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 19430 33200 19486 34000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 19982 33200 20038 34000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 20534 33200 20590 34000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5630 33200 5686 34000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 21086 33200 21142 34000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 21638 33200 21694 34000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 22190 33200 22246 34000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 22742 33200 22798 34000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 23294 33200 23350 34000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 23846 33200 23902 34000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 24398 33200 24454 34000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 24950 33200 25006 34000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 6182 33200 6238 34000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6734 33200 6790 34000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 7286 33200 7342 34000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 7838 33200 7894 34000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 8390 33200 8446 34000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 8942 33200 8998 34000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 9494 33200 9550 34000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4710 33200 4766 34000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 10230 33200 10286 34000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 10782 33200 10838 34000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 11334 33200 11390 34000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 11886 33200 11942 34000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 12438 33200 12494 34000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 12990 33200 13046 34000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 13542 33200 13598 34000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 14094 33200 14150 34000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 14646 33200 14702 34000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 15198 33200 15254 34000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5262 33200 5318 34000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 15750 33200 15806 34000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 16302 33200 16358 34000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 16854 33200 16910 34000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 17406 33200 17462 34000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 17958 33200 18014 34000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 18510 33200 18566 34000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 19062 33200 19118 34000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 19614 33200 19670 34000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 20166 33200 20222 34000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 20718 33200 20774 34000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 5814 33200 5870 34000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 21270 33200 21326 34000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 21822 33200 21878 34000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 22374 33200 22430 34000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 22926 33200 22982 34000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 23478 33200 23534 34000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 24030 33200 24086 34000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 24582 33200 24638 34000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 25134 33200 25190 34000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 6366 33200 6422 34000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 6918 33200 6974 34000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 7470 33200 7526 34000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 8022 33200 8078 34000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 8574 33200 8630 34000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 9126 33200 9182 34000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 9678 33200 9734 34000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4894 33200 4950 34000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 10414 33200 10470 34000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 10966 33200 11022 34000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 11518 33200 11574 34000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 12070 33200 12126 34000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 12622 33200 12678 34000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 13174 33200 13230 34000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 13726 33200 13782 34000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 14278 33200 14334 34000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 14830 33200 14886 34000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 15382 33200 15438 34000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5446 33200 5502 34000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 15934 33200 15990 34000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 16486 33200 16542 34000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 17038 33200 17094 34000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 17590 33200 17646 34000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 18142 33200 18198 34000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 18694 33200 18750 34000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 19246 33200 19302 34000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 19798 33200 19854 34000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 20350 33200 20406 34000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 20902 33200 20958 34000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 5998 33200 6054 34000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 21454 33200 21510 34000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 22006 33200 22062 34000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 22558 33200 22614 34000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 23110 33200 23166 34000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 23662 33200 23718 34000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 24214 33200 24270 34000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 24766 33200 24822 34000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 25318 33200 25374 34000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 6550 33200 6606 34000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 7102 33200 7158 34000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 7654 33200 7710 34000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 8206 33200 8262 34000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 8758 33200 8814 34000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 9310 33200 9366 34000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 9862 33200 9918 34000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4417 2128 4737 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 31600 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 34000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 495192
string GDS_FILE /home/runner/work/xls_workshop_tapeout_test_all_branch/xls_workshop_tapeout_test_all_branch/openlane/tiny_user_project/runs/22_12_16_09_52/results/signoff/tiny_user_project.magic.gds
string GDS_START 23768
<< end >>

